library IEEE;
use IEEE.STD_LOGIC_1164.all;

package InstructionMemory is


constant addr_max : integer := 103;
type IMtype is array (0 to addr_max) of std_logic_vector(31 downto 0);

constant IM : IMtype:= (X"03DEF026", X"03BDE826", X"039CE026", X"00000000", X"27DE0003", 
X"27BD0003", X"00000000", X"00000000", X"43DE000C", X"43BD000C", X"00000000", X"00000000", 
X"00000000", X"AFBEFFFC", X"AFBFFFF8", X"23DDFFF8", X"0C000005", X"00000000", X"AFA10000", 
X"0C000052", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", 
X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", X"3C020000", X"00000000", 
X"00000000", X"00000000", X"34420000", X"3C010000", X"00000000", X"00000000", X"00000000", 
X"34210004", X"00000000", X"00000000", X"00000000", X"8C420000", X"8C210000", X"00000000", 
X"00000000", X"00000000", X"0041D82A", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"08000010", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"3C1C0000", X"00000000", X"00000000", X"00000000", 
X"379C0001", X"0800000F", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"3C1C0000", X"00000000", X"00000000", X"00000000", X"379C0000", X"00000000", 
X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", 
X"00000000", X"03E00008", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"FFFFFFFF");


end InstructionMemory;
