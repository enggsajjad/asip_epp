library IEEE;
use IEEE.STD_LOGIC_1164.all;

package InstructionMemory is


constant addr_max : integer := 178;
type IMtype is array (0 to addr_max) of std_logic_vector(31 downto 0);

constant IM : IMtype:= (X"03DEF026", X"03BDE826", X"039CE026", X"00000000", X"27DE0003", 
X"27BD0003", X"00000000", X"00000000", X"43DE000C", X"43BD000C", X"00000000", X"00000000", 
X"00000000", X"AFBEFFFC", X"AFBFFFF8", X"23DDFFF8", X"0C000038", X"00000000", X"AFA10000", 
X"0C00009D", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", 
X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", X"0022D82B", X"00000000", 
X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", X"00000000", X"08000009", 
X"00000000", X"00000000", X"00000000", X"00201020", X"08000007", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"0040E020", X"00000000", X"00000000", 
X"00000000", X"08000004", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", 
X"03E00008", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"AFBEFFFC", X"AFBF0000", X"2FBE0004", X"2BBD000C", X"00000000", X"00000000", X"00000000", 
X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50008", X"00000000", X"00000000", 
X"3C010000", X"00000000", X"00000000", X"00000000", X"34210000", X"00000000", X"00000000", 
X"3C020000", X"00000000", X"00000000", X"00000000", X"34420004", X"3C040000", X"00000000", 
X"00000000", X"00000000", X"34840004", X"3C030000", X"00000000", X"00000000", X"00000000", 
X"34630000", X"00000000", X"00000000", X"00000000", X"AFC5FFFC", X"3C050000", X"00000000", 
X"00000000", X"00000000", X"34A50005", X"00000000", X"00000000", X"3C060000", X"00000000", 
X"00000000", X"00000000", X"34C60007", X"00000000", X"00000000", X"AC250000", X"00000000", 
X"00000000", X"00000000", X"AC460000", X"00000000", X"00000000", X"00000000", X"8C820000", 
X"8C610000", X"00000000", X"00000000", X"00000000", X"2BBD0008", X"00000000", X"00000000", 
X"00000000", X"0FFFFF83", X"00000000", X"00000000", X"00000000", X"23BD0008", X"00000000", 
X"00000000", X"00000000", X"8FC1FFFC", X"00000000", X"00000000", X"00000000", X"AC3C0000", 
X"08000004", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", X"03E00008", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"FFFFFFFF");


end InstructionMemory;
