library IEEE;
use IEEE.STD_LOGIC_1164.all;

package InstructionMemory is


constant addr_max : integer := 359;
type IMtype is array (0 to addr_max) of std_logic_vector(31 downto 0);

constant IM : IMtype:= (X"03DEF026", X"03BDE826", X"039CE026", X"00000000", X"3C1E000F", 
X"3C1D000F", X"00000000", X"00000000", X"37DEFFFC", X"37BDFFFC", X"00000000", X"00000000", 
X"00000000", X"AFBEFFFC", X"AFBFFFF8", X"23DDFFF8", X"0C000005", X"00000000", X"AFA10000", 
X"0C000152", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", 
X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", X"3C020000", X"00000000", 
X"00000000", X"00000000", X"3442FF00", X"3C010000", X"00000000", X"00000000", X"00000000", 
X"34210000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"3C030000", 
X"00000000", X"00000000", X"00000000", X"34630000", X"3C060000", X"00000000", X"00000000", 
X"00000000", X"34C60050", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840004", 
X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50004", X"00000000", X"00000000", 
X"00000000", X"00242018", X"00252818", X"3C070000", X"00000000", X"00000000", X"00000000", 
X"34E70004", X"3C080000", X"00000000", X"00000000", X"00000000", X"350800A0", X"00641820", 
X"00C52020", X"00273018", X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50004", 
X"8C630000", X"8C840000", X"01063020", X"3C070000", X"00000000", X"00000000", X"00000000", 
X"34E70000", X"00252818", X"C4641800", X"00000000", X"00000000", X"00000000", X"ACC30000", 
X"00E51820", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840004", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A500F0", X"00000000", X"00000000", X"8C630000", 
X"00242018", X"3C070000", X"00000000", X"00000000", X"00000000", X"34E70004", X"3C060000", 
X"00000000", X"00000000", X"00000000", X"34C60004", X"3C080000", X"00000000", X"00000000", 
X"00000000", X"35080004", X"00A42020", X"CC621A00", X"3C0A0000", X"00000000", X"00000000", 
X"00000000", X"354A0050", X"00273818", X"00000000", X"00000000", X"00000000", X"3C090000", 
X"00000000", X"00000000", X"00000000", X"35290000", X"00263018", X"AC830000", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50140", X"00284018", X"01472020", X"3C0B0000", 
X"00000000", X"00000000", X"00000000", X"356B0004", X"3C0C0000", X"00000000", X"00000000", 
X"00000000", X"358C0004", X"01261820", X"00A82820", X"8C840000", X"3C070000", X"00000000", 
X"00000000", X"00000000", X"34E70050", X"002C5018", X"3C060000", X"00000000", X"00000000", 
X"00000000", X"34C60000", X"002B4818", X"8C630000", X"00000000", X"00000000", X"00000000", 
X"C0641800", X"00000000", X"00000000", X"00000000", X"ACA30000", X"00EA2020", X"00C91820", 
X"00000000", X"00000000", X"00000000", X"8C840000", X"8C630000", X"00000000", X"00000000", 
X"00000000", X"0064D82A", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", 
X"00000000", X"00000000", X"08000030", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630000", X"3C040000", 
X"00000000", X"00000000", X"00000000", X"34840190", X"3C050000", X"00000000", X"00000000", 
X"00000000", X"34A50004", X"3C060000", X"00000000", X"00000000", X"00000000", X"34C60004", 
X"00000000", X"00000000", X"00000000", X"00252818", X"00263018", X"00000000", X"00000000", 
X"00000000", X"00651820", X"00862020", X"00000000", X"00000000", X"00000000", X"8C630000", 
X"00000000", X"00000000", X"00000000", X"AC830000", X"08000033", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", 
X"34630050", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840190", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50004", X"3C060000", X"00000000", X"00000000", 
X"00000000", X"34C60004", X"00000000", X"00000000", X"00000000", X"00252818", X"00263018", 
X"00000000", X"00000000", X"00000000", X"00651820", X"00862020", X"00000000", X"00000000", 
X"00000000", X"8C630000", X"00000000", X"00000000", X"00000000", X"AC830000", X"08000007", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"20210001", 
X"00000000", X"00000000", X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", 
X"34630014", X"00000000", X"00000000", X"00000000", X"0023D82A", X"00000000", X"00000000", 
X"00000000", X"1760FEEB", X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"3C1C0000", X"00000000", 
X"00000000", X"00000000", X"379C0000", X"00000000", X"00000000", X"00000000", X"08000004", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"8FDF0004", 
X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", X"03E00008", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"FFFFFFFF");


end InstructionMemory;
