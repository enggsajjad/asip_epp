library IEEE;
use IEEE.STD_LOGIC_1164.all;

package InstructionMemory is


constant addr_max : integer := 840;
type IMtype is array (0 to addr_max) of std_logic_vector(31 downto 0);

constant IM : IMtype:= (X"03DEF026", X"03BDE826", X"039CE026", X"00000000", X"27DE0003", 
X"27BD0003", X"00000000", X"00000000", X"43DE000C", X"43BD000C", X"00000000", X"00000000", 
X"00000000", X"AFBEFFFC", X"AFBFFFF8", X"23DDFFF8", X"0C00027C", X"00000000", X"AFA10000", 
X"0C000333", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", 
X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", X"40430008", X"3C020000", 
X"00000000", X"00000000", X"00000000", X"34420000", X"00000000", X"00000000", X"00000000", 
X"0061E026", X"00000000", X"00000000", X"00000000", X"33818000", X"00000000", X"00000000", 
X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630000", X"00000000", 
X"00000000", X"00000000", X"0023D82F", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"08000010", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"43810001", X"00000000", X"00000000", X"00000000", 
X"383C1021", X"0800000B", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"439C0001", X"00000000", X"00000000", X"00000000", X"20420001", X"00000000", 
X"00000000", X"00000000", X"3C010000", X"00000000", X"00000000", X"00000000", X"34210008", 
X"00000000", X"00000000", X"00000000", X"0041D82A", X"00000000", X"00000000", X"00000000", 
X"1760FFC5", X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", 
X"00000000", X"08000004", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", 
X"03E00008", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"AFBEFFFC", X"AFBF0000", X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", 
X"00202820", X"00000000", X"00000000", X"00000000", X"3C060000", X"00000000", X"00000000", 
X"00000000", X"34C60300", X"00000000", X"00000000", X"00000000", X"8CC10000", X"3C070000", 
X"00000000", X"00000000", X"00000000", X"34E70000", X"00000000", X"00000000", X"00000000", 
X"0027D82E", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", 
X"00000000", X"08000083", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"3C070000", X"00000000", X"00000000", X"00000000", X"34E70001", X"3C010000", 
X"00000000", X"00000000", X"00000000", X"34210000", X"00000000", X"00000000", X"00000000", 
X"ACC70000", X"08000062", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"40C60001", X"00000000", X"00000000", X"00000000", X"20E70001", X"00000000", 
X"00000000", X"00000000", X"3C080000", X"00000000", X"00000000", X"00000000", X"35080008", 
X"00000000", X"00000000", X"00000000", X"00E8D82A", X"00000000", X"00000000", X"00000000", 
X"17600184", X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", 
X"00000000", X"00204020", X"3C090000", X"00000000", X"00000000", X"00000000", X"35290100", 
X"3C070000", X"00000000", X"00000000", X"00000000", X"34E70404", X"00000000", X"00000000", 
X"00000000", X"302A000F", X"00205820", X"3C0C0000", X"00000000", X"00000000", X"00000000", 
X"358C0304", X"442D0004", X"00000000", X"00000000", X"00000000", X"20210001", X"00000000", 
X"00000000", X"00000000", X"00EA5020", X"00000000", X"00000000", X"41080001", X"00ED3820", 
X"00000000", X"00000000", X"00000000", X"01284020", X"00000000", X"00000000", X"00000000", 
X"A5060000", X"018B4820", X"00000000", X"00000000", X"00000000", X"81460000", X"80E70000", 
X"00000000", X"00000000", X"00000000", X"40C60004", X"00000000", X"00000000", X"00000000", 
X"00C73025", X"00000000", X"00000000", X"00000000", X"A1260000", X"00000000", X"00000000", 
X"00000000", X"703B00FF", X"00000000", X"00000000", X"00000000", X"14200129", X"00000000", 
X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", X"00000000", X"747B0000", 
X"00000000", X"00000000", X"00000000", X"14600008", X"00000000", X"00000000", X"00000000", 
X"08000011", X"00000000", X"00000000", X"00000000", X"00600820", X"00000000", X"00000000", 
X"00000000", X"40210008", X"00000000", X"00000000", X"00000000", X"00232825", X"0800003D", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"3C010000", 
X"00000000", X"00000000", X"00000000", X"34210000", X"00000000", X"00000000", X"00000000", 
X"0081D82A", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", 
X"00000000", X"08000026", X"00000000", X"00000000", X"00000000", X"30A300FF", X"3C010000", 
X"00000000", X"00000000", X"00000000", X"34210304", X"00000000", X"00000000", X"00000000", 
X"44A50008", X"00000000", X"00000000", X"00000000", X"00231820", X"00000000", X"00000000", 
X"00000000", X"80630000", X"00250820", X"00000000", X"00000000", X"00000000", X"80210000", 
X"00000000", X"00000000", X"00000000", X"40630008", X"00000000", X"00000000", X"00000000", 
X"00612825", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"3C010000", X"00000000", X"00000000", X"00000000", X"34210001", X"0800003B", X"00000000", 
X"00000000", X"00000000", X"3C060000", X"00000000", X"00000000", X"00000000", X"34C60000", 
X"00201820", X"44A70008", X"00000000", X"00000000", X"00000000", X"00C31820", X"00000000", 
X"00000000", X"00000000", X"80630000", X"00000000", X"00000000", X"00000000", X"00671826", 
X"00000000", X"00000000", X"00000000", X"30A500FF", X"00000000", X"00000000", X"00000000", 
X"3C060000", X"00000000", X"00000000", X"00000000", X"34C60100", X"20210001", X"00000000", 
X"00000000", X"00000000", X"40630001", X"00000000", X"00000000", X"00000000", X"00C31820", 
X"00000000", X"00000000", X"00000000", X"84630000", X"00000000", X"00000000", X"00000000", 
X"40A50008", X"00000000", X"00000000", X"00000000", X"00A32826", X"00000000", X"00000000", 
X"00000000", X"0022D82C", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", 
X"00000000", X"00000000", X"08000042", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630000", 
X"00000000", X"00000000", X"00000000", X"0083D82A", X"00000000", X"00000000", X"00000000", 
X"17600008", X"00000000", X"00000000", X"00000000", X"0BFFFFAA", X"00000000", X"00000000", 
X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630000", X"00203020", 
X"3C070000", X"00000000", X"00000000", X"00000000", X"34E70304", X"00000000", X"00000000", 
X"00000000", X"44A80008", X"00000000", X"00000000", X"00000000", X"00661820", X"00000000", 
X"00000000", X"00000000", X"80630000", X"00000000", X"00000000", X"00000000", X"00E31820", 
X"00000000", X"00000000", X"00000000", X"80630000", X"00000000", X"00000000", X"00000000", 
X"00681826", X"0BFFFF99", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"3C010000", X"00000000", X"00000000", X"00000000", X"34210000", X"00000000", 
X"00000000", X"00000000", X"0081D82D", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"08000009", X"00000000", X"00000000", X"00000000", 
X"00A0E020", X"08000026", X"00000000", X"00000000", X"00000000", X"30A200FF", X"3C010000", 
X"00000000", X"00000000", X"00000000", X"34210304", X"00000000", X"00000000", X"00000000", 
X"44A30008", X"00000000", X"00000000", X"00000000", X"00221020", X"00000000", X"00000000", 
X"00000000", X"80420000", X"00230820", X"00000000", X"00000000", X"00000000", X"80210000", 
X"00000000", X"00000000", X"00000000", X"40420008", X"00000000", X"00000000", X"00000000", 
X"0041E025", X"00000000", X"00000000", X"00000000", X"08000038", X"00000000", X"00000000", 
X"00000000", X"00203020", X"00000000", X"00000000", X"00000000", X"3C070000", X"00000000", 
X"00000000", X"00000000", X"34E70000", X"00000000", X"00000000", X"00000000", X"40C60008", 
X"00000000", X"00000000", X"00000000", X"30C88000", X"00000000", X"00000000", X"00000000", 
X"3C090000", X"00000000", X"00000000", X"00000000", X"35290000", X"00000000", X"00000000", 
X"00000000", X"0109D82F", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", 
X"00000000", X"00000000", X"0BFFFE51", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"40C60001", X"00000000", X"00000000", X"00000000", X"38C61021", 
X"0BFFFE4C", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", X"03E00008", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", 
X"AFBF0000", X"2FBE0004", X"2BBD0014", X"00000000", X"00000000", X"00000000", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50000", X"00000000", X"00000000", X"3C010000", 
X"00000000", X"00000000", X"00000000", X"34210414", X"00000000", X"00000000", X"00000000", 
X"3C070000", X"00000000", X"00000000", X"00000000", X"34E70029", X"00000000", X"00000000", 
X"3C060000", X"00000000", X"00000000", X"00000000", X"34C60000", X"AFC1FFFC", X"00A72820", 
X"3C040000", X"00000000", X"00000000", X"00000000", X"34840001", X"3C030000", X"00000000", 
X"00000000", X"00000000", X"34630000", X"3C020000", X"00000000", X"00000000", X"00000000", 
X"34420028", X"3C010000", X"00000000", X"00000000", X"00000000", X"34210000", X"AFC5FFF8", 
X"A0A60000", X"00000000", X"00000000", X"00000000", X"2BBD0008", X"00000000", X"00000000", 
X"00000000", X"0FFFFDB0", X"00000000", X"00000000", X"00000000", X"23BD0008", X"00000000", 
X"00000000", X"00000000", X"8FC1FFFC", X"00000000", X"00000000", X"3C040000", X"00000000", 
X"00000000", X"00000000", X"34840416", X"00000000", X"00000000", X"A43C0000", X"00000000", 
X"00000000", X"00000000", X"84220000", X"00000000", X"00000000", X"00000000", X"00400820", 
X"44430008", X"304200FF", X"00000000", X"00000000", X"00000000", X"20630001", X"20450001", 
X"8FC2FFF8", X"00000000", X"00000000", X"00000000", X"00403820", X"A0430000", X"00000000", 
X"00000000", X"00000000", X"3C060000", X"00000000", X"00000000", X"00000000", X"34C60001", 
X"AFC4FFF4", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840001", X"00000000", 
X"00000000", X"00E63020", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630000", 
X"3C020000", X"00000000", X"00000000", X"00000000", X"3442002A", X"00000000", X"00000000", 
X"A0C50000", X"00000000", X"00000000", X"00000000", X"2BBD0008", X"00000000", X"00000000", 
X"00000000", X"0FFFFD63", X"00000000", X"00000000", X"00000000", X"23BD0008", X"00000000", 
X"00000000", X"00000000", X"8FC1FFF4", X"00000000", X"00000000", X"00000000", X"A43C0000", 
X"00000000", X"00000000", X"00000000", X"3C1C0000", X"00000000", X"00000000", X"00000000", 
X"379C0000", X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"8FDF0004", X"27DD0004", X"8FDE0000", 
X"00000000", X"00000000", X"00000000", X"03E00008", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"FFFFFFFF");


end InstructionMemory;
