library IEEE;
use IEEE.STD_LOGIC_1164.all;

package InstructionMemory is


constant addr_max : integer := 1051;
type IMtype is array (0 to addr_max) of std_logic_vector(31 downto 0);

constant IM : IMtype:= (X"03DEF026", X"03BDE826", X"039CE026", X"00000000", X"27DE0003", 
X"27BD0003", X"00000000", X"00000000", X"43DE000C", X"43BD000C", X"00000000", X"00000000", 
X"00000000", X"AFBEFFFC", X"AFBFFFF8", X"23DDFFF8", X"0C000268", X"00000000", X"AFA10000", 
X"0C000406", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", 
X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", X"40430008", X"3C020000", 
X"00000000", X"00000000", X"00000000", X"34420008", X"00000000", X"00000000", X"00000000", 
X"0061E026", X"00000000", X"00000000", X"00000000", X"33818000", X"00000000", X"00000000", 
X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630000", X"00000000", 
X"00000000", X"00000000", X"0023D82F", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"08000090", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"43810001", X"00000000", X"00000000", X"00000000", 
X"38211021", X"00000000", X"00000000", X"00000000", X"30238000", X"00000000", X"00000000", 
X"00000000", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840000", X"00000000", 
X"00000000", X"00000000", X"0064D82F", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"08000075", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"40210001", X"00000000", X"00000000", X"00000000", 
X"38211021", X"00000000", X"00000000", X"00000000", X"30238000", X"00000000", X"00000000", 
X"00000000", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840000", X"00000000", 
X"00000000", X"00000000", X"0064D82F", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"0800005A", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"40210001", X"00000000", X"00000000", X"00000000", 
X"38211021", X"00000000", X"00000000", X"00000000", X"30238000", X"00000000", X"00000000", 
X"00000000", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840000", X"00000000", 
X"00000000", X"00000000", X"0064D82F", X"00000000", X"00000000", X"00000000", X"17600008", 
X"00000000", X"00000000", X"00000000", X"0800003F", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"40210001", X"00000000", X"00000000", X"00000000", 
X"383C1021", X"00000000", X"00000000", X"00000000", X"2042FFFC", X"00000000", X"00000000", 
X"00000000", X"3C010000", X"00000000", X"00000000", X"00000000", X"34210000", X"00000000", 
X"00000000", X"00000000", X"0041D82B", X"00000000", X"00000000", X"00000000", X"1760FF64", 
X"00000000", X"00000000", X"00000000", X"08000024", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"43810001", X"0BFFFF7B", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40210001", X"0BFFFF96", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"40210001", X"0BFFFFB1", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"403C0001", 
X"0BFFFFCC", X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"8FDF0004", X"27DD0004", X"8FDE0000", 
X"00000000", X"00000000", X"00000000", X"03E00008", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", X"2FBE0004", X"2BBD0008", 
X"00000000", X"00000000", X"00000000", X"3C020000", X"00000000", X"00000000", X"00000000", 
X"3442022C", X"00000000", X"00000000", X"00000000", X"8C410000", X"3C030000", X"00000000", 
X"00000000", X"00000000", X"34630000", X"00000000", X"00000000", X"00000000", X"0023D82E", 
X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", X"00000000", 
X"08000064", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"3C030000", X"00000000", X"00000000", X"00000000", X"34630001", X"3C010000", X"00000000", 
X"00000000", X"00000000", X"34210000", X"00000000", X"00000000", X"00000000", X"AC430000", 
X"08000043", X"00000000", X"00000000", X"00000000", X"00202020", X"3C050000", X"00000000", 
X"00000000", X"00000000", X"34A5002A", X"3C030000", X"00000000", X"00000000", X"00000000", 
X"34630330", X"00000000", X"00000000", X"00000000", X"3026000F", X"00203820", X"3C080000", 
X"00000000", X"00000000", X"00000000", X"35080230", X"44290004", X"00000000", X"00000000", 
X"00000000", X"20210001", X"00000000", X"00000000", X"00000000", X"00663020", X"00000000", 
X"00000000", X"40840001", X"00691820", X"00000000", X"00000000", X"00000000", X"00A42020", 
X"00000000", X"00000000", X"00000000", X"A4820000", X"01072820", X"00000000", X"00000000", 
X"00000000", X"80C20000", X"80630000", X"00000000", X"00000000", X"00000000", X"40420004", 
X"00000000", X"00000000", X"00000000", X"00431025", X"00000000", X"00000000", X"00000000", 
X"A0A20000", X"00000000", X"00000000", X"00000000", X"703B0005", X"00000000", X"00000000", 
X"00000000", X"17600017", X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"3C1C0000", X"00000000", 
X"00000000", X"00000000", X"379C0000", X"00000000", X"00000000", X"00000000", X"080000D8", 
X"00000000", X"00000000", X"00000000", X"00201020", X"00000000", X"00000000", X"00000000", 
X"3C030000", X"00000000", X"00000000", X"00000000", X"34630008", X"00000000", X"00000000", 
X"00000000", X"40420008", X"00000000", X"00000000", X"00000000", X"30448000", X"00000000", 
X"00000000", X"00000000", X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50000", 
X"00000000", X"00000000", X"00000000", X"0085D82F", X"00000000", X"00000000", X"00000000", 
X"17600008", X"00000000", X"00000000", X"00000000", X"08000090", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"00000000", X"00000000", 
X"00000000", X"38421021", X"00000000", X"00000000", X"00000000", X"30448000", X"00000000", 
X"00000000", X"00000000", X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50000", 
X"00000000", X"00000000", X"00000000", X"0085D82F", X"00000000", X"00000000", X"00000000", 
X"17600008", X"00000000", X"00000000", X"00000000", X"08000075", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"00000000", X"00000000", 
X"00000000", X"38421021", X"00000000", X"00000000", X"00000000", X"30448000", X"00000000", 
X"00000000", X"00000000", X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50000", 
X"00000000", X"00000000", X"00000000", X"0085D82F", X"00000000", X"00000000", X"00000000", 
X"17600008", X"00000000", X"00000000", X"00000000", X"0800005A", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"00000000", X"00000000", 
X"00000000", X"38421021", X"00000000", X"00000000", X"00000000", X"30448000", X"00000000", 
X"00000000", X"00000000", X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50000", 
X"00000000", X"00000000", X"00000000", X"0085D82F", X"00000000", X"00000000", X"00000000", 
X"17600008", X"00000000", X"00000000", X"00000000", X"0800003F", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"00000000", X"00000000", 
X"00000000", X"38421021", X"00000000", X"00000000", X"00000000", X"2063FFFC", X"00000000", 
X"00000000", X"00000000", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840000", 
X"00000000", X"00000000", X"00000000", X"0064D82B", X"00000000", X"00000000", X"00000000", 
X"1760FF64", X"00000000", X"00000000", X"00000000", X"0BFFFEF6", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"0BFFFF7B", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"0BFFFF96", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", 
X"0BFFFFB1", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"40420001", X"0BFFFFCC", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", 
X"03E00008", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"AFBEFFFC", X"AFBF0000", X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", 
X"3C010000", X"00000000", X"00000000", X"00000000", X"34210000", X"00000000", X"00000000", 
X"3C020000", X"00000000", X"00000000", X"00000000", X"3442022C", X"00000000", X"00000000", 
X"00000000", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630029", X"00000000", 
X"00000000", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840000", X"00000000", 
X"00000000", X"00230820", X"3C050000", X"00000000", X"00000000", X"00000000", X"34A50000", 
X"00000000", X"00000000", X"00000000", X"A0240000", X"00000000", X"00000000", X"00000000", 
X"8C410000", X"00000000", X"00000000", X"00000000", X"0025D82E", X"00000000", X"00000000", 
X"00000000", X"17600008", X"00000000", X"00000000", X"00000000", X"08000064", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"3C030000", X"00000000", 
X"00000000", X"00000000", X"34630001", X"3C010000", X"00000000", X"00000000", X"00000000", 
X"34210000", X"00000000", X"00000000", X"00000000", X"AC430000", X"08000043", X"00000000", 
X"00000000", X"00000000", X"00202020", X"3C050000", X"00000000", X"00000000", X"00000000", 
X"34A5002A", X"3C030000", X"00000000", X"00000000", X"00000000", X"34630330", X"00000000", 
X"00000000", X"00000000", X"3026000F", X"00203820", X"3C080000", X"00000000", X"00000000", 
X"00000000", X"35080230", X"44290004", X"00000000", X"00000000", X"00000000", X"20210001", 
X"00000000", X"00000000", X"00000000", X"00663020", X"00000000", X"00000000", X"40840001", 
X"00691820", X"00000000", X"00000000", X"00000000", X"00A42020", X"00000000", X"00000000", 
X"00000000", X"A4820000", X"01072820", X"00000000", X"00000000", X"00000000", X"80C20000", 
X"80630000", X"00000000", X"00000000", X"00000000", X"40420004", X"00000000", X"00000000", 
X"00000000", X"00431025", X"00000000", X"00000000", X"00000000", X"A0A20000", X"00000000", 
X"00000000", X"00000000", X"703B0005", X"00000000", X"00000000", X"00000000", X"17600024", 
X"00000000", X"00000000", X"00000000", X"08000004", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"3C010000", X"00000000", X"00000000", X"00000000", X"34210340", 
X"00000000", X"00000000", X"00000000", X"3C020000", X"00000000", X"00000000", X"00000000", 
X"34420000", X"3C1C0000", X"00000000", X"00000000", X"00000000", X"379C0000", X"00000000", 
X"00000000", X"00000000", X"A4220000", X"080000D8", X"00000000", X"00000000", X"00000000", 
X"00201020", X"00000000", X"00000000", X"00000000", X"3C030000", X"00000000", X"00000000", 
X"00000000", X"34630008", X"00000000", X"00000000", X"00000000", X"40420008", X"00000000", 
X"00000000", X"00000000", X"30448000", X"00000000", X"00000000", X"00000000", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50000", X"00000000", X"00000000", X"00000000", 
X"0085D82F", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", 
X"00000000", X"08000090", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"40420001", X"00000000", X"00000000", X"00000000", X"38421021", X"00000000", 
X"00000000", X"00000000", X"30448000", X"00000000", X"00000000", X"00000000", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50000", X"00000000", X"00000000", X"00000000", 
X"0085D82F", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", 
X"00000000", X"08000075", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"40420001", X"00000000", X"00000000", X"00000000", X"38421021", X"00000000", 
X"00000000", X"00000000", X"30448000", X"00000000", X"00000000", X"00000000", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50000", X"00000000", X"00000000", X"00000000", 
X"0085D82F", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", 
X"00000000", X"0800005A", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"40420001", X"00000000", X"00000000", X"00000000", X"38421021", X"00000000", 
X"00000000", X"00000000", X"30448000", X"00000000", X"00000000", X"00000000", X"3C050000", 
X"00000000", X"00000000", X"00000000", X"34A50000", X"00000000", X"00000000", X"00000000", 
X"0085D82F", X"00000000", X"00000000", X"00000000", X"17600008", X"00000000", X"00000000", 
X"00000000", X"0800003F", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"40420001", X"00000000", X"00000000", X"00000000", X"38421021", X"00000000", 
X"00000000", X"00000000", X"2063FFFC", X"00000000", X"00000000", X"00000000", X"3C040000", 
X"00000000", X"00000000", X"00000000", X"34840000", X"00000000", X"00000000", X"00000000", 
X"0064D82B", X"00000000", X"00000000", X"00000000", X"1760FF64", X"00000000", X"00000000", 
X"00000000", X"0BFFFEE9", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"40420001", X"0BFFFF7B", X"00000000", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"40420001", X"0BFFFF96", X"00000000", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"40420001", X"0BFFFFB1", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"40420001", X"0BFFFFCC", X"00000000", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"8FDF0004", X"27DD0004", 
X"8FDE0000", X"00000000", X"00000000", X"00000000", X"03E00008", X"00000000", X"00000000", 
X"00000000", X"00000000", X"00000000", X"FFFFFFFF");


end InstructionMemory;
