library IEEE;
use IEEE.STD_LOGIC_1164.all;

package InstructionMemory is


constant addr_max : integer := 150;
type IMtype is array (0 to addr_max) of std_logic_vector(31 downto 0);

constant IM : IMtype:= (X"03DEF026", X"03BDE826", X"039CE026", X"00000000", X"27DE0003", 
X"27BD0003", X"00000000", X"00000000", X"43DE000C", X"43BD000C", X"00000000", X"00000000", 
X"00000000", X"AFBEFFFC", X"AFBFFFF8", X"23DDFFF8", X"0C000005", X"00000000", X"AFA10000", 
X"0C000081", X"00000000", X"00000000", X"00000000", X"00000000", X"AFBEFFFC", X"AFBF0000", 
X"2FBE0004", X"2BBD0008", X"00000000", X"00000000", X"00000000", X"3C010000", X"00000000", 
X"00000000", X"00000000", X"34210000", X"00000000", X"00000000", X"3C020000", X"00000000", 
X"00000000", X"00000000", X"34420004", X"00000000", X"00000000", X"3C030000", X"00000000", 
X"00000000", X"00000000", X"34630008", X"3C050000", X"00000000", X"00000000", X"00000000", 
X"34A50000", X"3C040000", X"00000000", X"00000000", X"00000000", X"34840004", X"3C060000", 
X"00000000", X"00000000", X"00000000", X"34C60008", X"3C070000", X"00000000", X"00000000", 
X"00000000", X"34E70008", X"3C080000", X"00000000", X"00000000", X"00000000", X"35080008", 
X"00000000", X"00000000", X"00000000", X"3C090000", X"00000000", X"00000000", X"00000000", 
X"35290003", X"00000000", X"00000000", X"3C0A0000", X"00000000", X"00000000", X"00000000", 
X"354A0005", X"00000000", X"00000000", X"AC290000", X"3C0B0000", X"00000000", X"00000000", 
X"00000000", X"356B0007", X"00000000", X"00000000", X"00000000", X"AC4A0000", X"00000000", 
X"00000000", X"00000000", X"AC6B0000", X"00000000", X"00000000", X"00000000", X"8CA10000", 
X"8C820000", X"8CC30000", X"00000000", X"00000000", X"00000000", X"00220818", X"00000000", 
X"00000000", X"00000000", X"00610820", X"00000000", X"00000000", X"00000000", X"ACE10000", 
X"00000000", X"00000000", X"00000000", X"8D1C0000", X"00000000", X"00000000", X"00000000", 
X"08000004", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", 
X"8FDF0004", X"27DD0004", X"8FDE0000", X"00000000", X"00000000", X"00000000", X"03E00008", 
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"FFFFFFFF");


end InstructionMemory;
