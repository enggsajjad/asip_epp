--   int_port : internal port
--   ext_port : external port

-- Comment :

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.numeric_std.all;

entity fhm_rotator_w32 is
  port (
data_in   : in  std_logic_vector(31 downto 0);
direction : in  std_logic;
amount    : in  std_logic_vector(7 downto 0);
data_out  : out std_logic_vector(31 downto 0)
        );
end fhm_rotator_w32;

architecture logic of fhm_rotator_w32 is

begin
  process (data_in, amount, direction)
variable a    : integer;
variable res : std_logic_vector(31 downto 0);
begin
     a := TO_INTEGER(UNSIGNED(amount));
     if (a > 0 and a < 32) then
          case direction is
          when '0' => -- rotate left
               res(31 - a downto 0) :=
                    data_in(31 downto a);
               res(31 downto 32 - a) :=
                    data_in(a - 1 downto 0);
          when others => -- not reached
               res := (others => 'X');
          end case;
     else
          res := (others => 'X');
     end if;
     data_out <= res;
end process;

end logic;


-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
